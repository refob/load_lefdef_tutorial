VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X1 0 0 ;
  SIZE 3.2 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.3 0.6 4.1 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.3 4.9 1.7 5.7 ;
        RECT 1 5.3 1.7 5.7 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.5 -0.3 1.9 2.6 ;
        RECT -0.2 -0.3 3.4 0.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6 6.3 3 6.7 ;
        RECT 2.6 7.4 3 9.4 ;
        RECT 2.7 1.6 3 9.4 ;
        RECT 2.3 0.6 2.7 1.9 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 7.4 0.6 10.3 ;
        RECT -0.2 9.7 3.4 10.3 ;
        RECT 1.8 7.4 2.2 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.2 0.6 0.6 2.6 ;
      RECT 0.3 2.6 1.2 2.9 ;
      RECT 0.9 2.6 1.2 3.3 ;
      RECT 2 2.9 2.4 3.3 ;
      RECT 0.9 3 2.4 3.3 ;
      RECT 2 2.9 2.3 7.1 ;
      RECT 1.1 6.8 2.3 7.1 ;
      RECT 1.1 6.8 1.4 9.4 ;
      RECT 1 7.4 1.4 9.4 ;
  END
END AND2X1

MACRO AND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X2 0 0 ;
  SIZE 3.2 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.3 0.6 4.1 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.1 3.6 1.4 4.7 ;
        RECT 1.2 3.5 1.6 3.9 ;
        RECT 1 4.3 1.4 4.7 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.5 -0.3 1.9 2.5 ;
        RECT -0.2 -0.3 3.4 0.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6 4.3 3 4.7 ;
        RECT 2.6 5.4 3 9.4 ;
        RECT 2.7 2.1 3 9.4 ;
        RECT 2.3 0.6 2.7 2.6 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 7.4 0.6 10.3 ;
        RECT -0.2 9.7 3.4 10.3 ;
        RECT 1.8 5.6 2.2 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.2 0.6 0.6 2.6 ;
      RECT 0.3 0.6 0.6 3 ;
      RECT 0.3 2.7 1.2 3 ;
      RECT 0.9 2.9 2.4 3.2 ;
      RECT 2 2.9 2.4 3.3 ;
      RECT 2 2.9 2.3 5.3 ;
      RECT 1.1 5 2.3 5.3 ;
      RECT 1.1 5 1.4 9.4 ;
      RECT 1 7.4 1.4 9.4 ;
  END
END AND2X2

MACRO AOI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X1 0 0 ;
  SIZE 3.2 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 4.3 0.6 4.7 ;
        RECT 0.6 4.4 1 4.9 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 3.3 1.4 4.1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.5 1.9 2.9 2.3 ;
        RECT 2.6 2.3 3 2.7 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.5 -0.3 0.9 2.6 ;
        RECT -0.2 -0.3 3.4 0.3 ;
        RECT 2.6 -0.3 3 1.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 0.6 2.1 4.7 ;
        RECT 2.6 5.4 3 9.4 ;
        RECT 1.8 4.4 3 4.7 ;
        RECT 2.6 4.3 3 4.7 ;
        RECT 2.6 4.3 2.9 9.4 ;
        RECT 1.8 0.6 2.2 2.6 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 6 1.4 10.3 ;
        RECT -0.2 9.7 3.4 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.2 5.4 2.2 5.7 ;
      RECT 0.2 5.4 0.6 9.4 ;
      RECT 1.8 5.4 2.2 9.4 ;
  END
END AOI21X1

MACRO AOI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X1 0 0 ;
  SIZE 4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 4.3 0.6 4.7 ;
        RECT 0.6 4.4 1 4.9 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 3.3 1.4 4.1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.4 4.3 3.8 5.1 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6 3.3 2.9 4.3 ;
        RECT 2.6 3.3 3 3.7 ;
        RECT 2.5 3.9 2.9 4.3 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.4 -0.3 0.8 2.6 ;
        RECT -0.2 -0.3 4.2 0.3 ;
        RECT 3.4 -0.3 3.8 2.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 4.3 2.2 4.7 ;
        RECT 2.6 5.4 3 8.8 ;
        RECT 2.6 4.8 2.9 8.8 ;
        RECT 1.9 4.8 2.9 5.1 ;
        RECT 1.7 0.6 2.5 2.6 ;
        RECT 1.9 0.6 2.2 5.1 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 6 1.4 10.3 ;
        RECT -0.2 9.7 4.2 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.2 5.4 2.2 5.7 ;
      RECT 1.8 5.4 2.2 9.4 ;
      RECT 0.2 5.4 0.6 9.4 ;
      RECT 3.4 5.4 3.8 9.4 ;
      RECT 1.8 9.1 3.8 9.4 ;
  END
END AOI22X1

MACRO BUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2 0 0 ;
  SIZE 2.4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.9 0.6 4.7 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 2.6 ;
        RECT -0.2 -0.3 2.6 0.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 0.6 2.2 4.3 ;
        RECT 1.8 5.4 2.2 9.4 ;
        RECT 1.9 0.6 2.2 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 6 1.4 10.3 ;
        RECT -0.2 9.7 2.6 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.2 0.6 0.6 3.2 ;
      RECT 0.2 2.9 1.3 3.2 ;
      RECT 1 4.7 1.6 5.1 ;
      RECT 1 2.9 1.3 5.7 ;
      RECT 0.2 5.4 1.3 5.7 ;
      RECT 0.2 5.4 0.6 9.4 ;
  END
END BUFX2

MACRO BUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX4 0 0 ;
  SIZE 3.2 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3 3.9 0.7 4.7 ;
        RECT 0.2 4.3 0.7 4.7 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 2.6 ;
        RECT -0.2 -0.3 3.4 0.3 ;
        RECT 2.6 -0.3 3 2.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 0.6 2.2 2.6 ;
        RECT 2 2.3 2.3 5.9 ;
        RECT 1.8 5.4 2.2 9.4 ;
        RECT 1.8 3.3 2.3 3.7 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 6 1.4 10.3 ;
        RECT -0.2 9.7 3.4 10.3 ;
        RECT 2.6 5.4 3 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.2 0.6 0.6 3.2 ;
      RECT 0.2 2.9 1.5 3.2 ;
      RECT 1.2 4 1.7 4.4 ;
      RECT 1.2 2.9 1.5 5.7 ;
      RECT 0.2 5.4 1.5 5.7 ;
      RECT 0.2 5.4 0.6 9.4 ;
  END
END BUFX4

MACRO CLKBUF1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF1 0 0 ;
  SIZE 7.2 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.3 0.6 4 ;
        RECT 0.2 3.6 1.1 4 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 2.6 ;
        RECT -0.2 -0.3 7.4 0.3 ;
        RECT 6.6 -0.3 7 2.6 ;
        RECT 5 -0.3 5.4 2.6 ;
        RECT 3.4 -0.3 3.8 2.6 ;
        RECT 1.8 -0.3 2.2 2.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.8 0.6 6.2 3.3 ;
        RECT 5.8 4.7 7 5.1 ;
        RECT 6.6 2.9 7 5.1 ;
        RECT 5.8 2.9 7 3.3 ;
        RECT 5.8 4.7 6.2 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 7.4 10.3 ;
        RECT 6.6 5.4 7 10.3 ;
        RECT 5 5.4 5.4 10.3 ;
        RECT 3.4 5.4 3.8 10.3 ;
        RECT 1.8 5.4 2.2 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 1 0.6 1.4 3.3 ;
      RECT 1 2.9 1.9 3.3 ;
      RECT 1.5 3.6 2.8 4 ;
      RECT 1.5 2.9 1.9 5.1 ;
      RECT 1 4.7 1.9 5.1 ;
      RECT 1 4.7 1.4 9.4 ;
      RECT 2.6 0.6 3 3.3 ;
      RECT 2.6 2.9 3.7 3.3 ;
      RECT 3.3 3.6 4.5 4 ;
      RECT 3.3 2.9 3.7 5.1 ;
      RECT 2.6 4.7 3.7 5.1 ;
      RECT 2.6 4.7 3 9.4 ;
      RECT 4.2 0.6 4.6 3.3 ;
      RECT 4.2 2.9 5.3 3.3 ;
      RECT 4.9 3.6 6.2 4 ;
      RECT 4.9 2.9 5.3 5.1 ;
      RECT 4.2 4.7 5.3 5.1 ;
      RECT 4.2 4.7 4.6 9.4 ;
  END
END CLKBUF1

MACRO CLKBUF2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF2 0 0 ;
  SIZE 10.4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.3 0.6 4 ;
        RECT 0.2 3.6 1.1 4 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 2.6 ;
        RECT -0.2 -0.3 10.6 0.3 ;
        RECT 9.8 -0.3 10.2 2.6 ;
        RECT 8.2 -0.3 8.6 2.6 ;
        RECT 6.6 -0.3 7 2.6 ;
        RECT 5 -0.3 5.4 2.6 ;
        RECT 3.4 -0.3 3.8 2.6 ;
        RECT 1.8 -0.3 2.2 2.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9 0.6 9.4 3.3 ;
        RECT 9 4.7 10.2 5.1 ;
        RECT 9.8 2.9 10.2 5.1 ;
        RECT 9 2.9 10.2 3.3 ;
        RECT 9 4.7 9.4 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 10.6 10.3 ;
        RECT 9.8 5.4 10.2 10.3 ;
        RECT 8.2 5.4 8.6 10.3 ;
        RECT 6.6 5.4 7 10.3 ;
        RECT 5 5.4 5.4 10.3 ;
        RECT 3.4 5.4 3.8 10.3 ;
        RECT 1.8 5.4 2.2 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 1 0.6 1.4 3.3 ;
      RECT 1 2.9 1.9 3.3 ;
      RECT 1.5 3.6 2.8 4 ;
      RECT 1.5 2.9 1.9 5.1 ;
      RECT 1 4.7 1.9 5.1 ;
      RECT 1 4.7 1.4 9.4 ;
      RECT 2.6 0.6 3 3.3 ;
      RECT 2.6 2.9 3.7 3.3 ;
      RECT 3.3 3.6 4.5 4 ;
      RECT 3.3 2.9 3.7 5.1 ;
      RECT 2.6 4.7 3.7 5.1 ;
      RECT 2.6 4.7 3 9.4 ;
      RECT 4.2 0.6 4.6 3.3 ;
      RECT 4.2 2.9 5.3 3.3 ;
      RECT 4.9 3.6 6.2 4 ;
      RECT 4.9 2.9 5.3 5.1 ;
      RECT 4.2 4.7 5.3 5.1 ;
      RECT 4.2 4.7 4.6 9.4 ;
      RECT 5.8 0.6 6.2 3.3 ;
      RECT 5.8 2.9 7 3.3 ;
      RECT 6.6 3.6 7.5 4 ;
      RECT 6.6 2.9 7 5.1 ;
      RECT 5.8 4.7 7 5.1 ;
      RECT 5.8 4.7 6.2 9.4 ;
      RECT 7.4 0.6 7.8 3.3 ;
      RECT 7.4 2.9 8.3 3.3 ;
      RECT 7.9 3.6 9.2 4 ;
      RECT 7.9 2.9 8.3 5.1 ;
      RECT 7.4 4.7 8.3 5.1 ;
      RECT 7.4 4.7 7.8 9.4 ;
  END
END CLKBUF2

MACRO CLKBUF3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF3 0 0 ;
  SIZE 13.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.3 0.6 4 ;
        RECT 0.2 3.6 1.1 4 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 2.6 ;
        RECT -0.2 -0.3 13.8 0.3 ;
        RECT 13 -0.3 13.4 2.6 ;
        RECT 11.4 -0.3 11.8 2.6 ;
        RECT 9.8 -0.3 10.2 2.6 ;
        RECT 8.2 -0.3 8.6 2.6 ;
        RECT 6.6 -0.3 7 2.6 ;
        RECT 5 -0.3 5.4 2.6 ;
        RECT 3.4 -0.3 3.8 2.6 ;
        RECT 1.8 -0.3 2.2 2.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.2 0.6 12.6 3.3 ;
        RECT 12.2 4.7 13.4 5.1 ;
        RECT 13 2.9 13.4 5.1 ;
        RECT 12.2 2.9 13.4 3.3 ;
        RECT 12.2 4.7 12.6 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 13.8 10.3 ;
        RECT 13 5.4 13.4 10.3 ;
        RECT 11.4 5.4 11.8 10.3 ;
        RECT 9.8 5.4 10.2 10.3 ;
        RECT 8.2 5.4 8.6 10.3 ;
        RECT 6.6 5.4 7 10.3 ;
        RECT 5 5.4 5.4 10.3 ;
        RECT 3.4 5.4 3.8 10.3 ;
        RECT 1.8 5.4 2.2 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 1 0.6 1.4 3.3 ;
      RECT 1 2.9 1.9 3.3 ;
      RECT 1.5 3.6 2.8 4 ;
      RECT 1.5 2.9 1.9 5.1 ;
      RECT 1 4.7 1.9 5.1 ;
      RECT 1 4.7 1.4 9.4 ;
      RECT 2.6 0.6 3 3.3 ;
      RECT 2.6 2.9 3.7 3.3 ;
      RECT 3.3 3.6 4.5 4 ;
      RECT 3.3 2.9 3.7 5.1 ;
      RECT 2.6 4.7 3.7 5.1 ;
      RECT 2.6 4.7 3 9.4 ;
      RECT 4.2 0.6 4.6 3.3 ;
      RECT 4.2 2.9 5.3 3.3 ;
      RECT 4.9 3.6 6.2 4 ;
      RECT 4.9 2.9 5.3 5.1 ;
      RECT 4.2 4.7 5.3 5.1 ;
      RECT 4.2 4.7 4.6 9.4 ;
      RECT 5.8 0.6 6.2 3.3 ;
      RECT 5.8 2.9 7 3.3 ;
      RECT 6.6 3.6 7.5 4 ;
      RECT 6.6 2.9 7 5.1 ;
      RECT 5.8 4.7 7 5.1 ;
      RECT 5.8 4.7 6.2 9.4 ;
      RECT 7.4 0.6 7.8 3.3 ;
      RECT 7.4 2.9 8.3 3.3 ;
      RECT 7.9 3.6 9.2 4 ;
      RECT 7.9 2.9 8.3 5.1 ;
      RECT 7.4 4.7 8.3 5.1 ;
      RECT 7.4 4.7 7.8 9.4 ;
      RECT 9 0.6 9.4 3.3 ;
      RECT 9 2.9 10.1 3.3 ;
      RECT 9.7 3.6 10.9 4 ;
      RECT 9.7 2.9 10.1 5.1 ;
      RECT 9 4.7 10.1 5.1 ;
      RECT 9 4.7 9.4 9.4 ;
      RECT 10.6 0.6 11 3.3 ;
      RECT 10.6 2.9 11.7 3.3 ;
      RECT 11.3 3.6 12.6 4 ;
      RECT 11.3 2.9 11.7 5.1 ;
      RECT 10.6 4.7 11.7 5.1 ;
      RECT 10.6 4.7 11 9.4 ;
  END
END CLKBUF3

MACRO DFFNEGX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNEGX1 0 0 ;
  SIZE 9.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.3 4.7 7.7 5.1 ;
        RECT 9 0.6 9.4 9.4 ;
        RECT 7.3 4.8 9.4 5.1 ;
        RECT 7.5 2.8 9.4 3.1 ;
        RECT 7.5 2.7 7.9 3.1 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal2 ;
        RECT 2.6 3.4 3 6.7 ;
      LAYER via ;
        RECT 2.7 6.4 2.9 6.6 ;
        RECT 2.7 3.5 2.9 3.7 ;
      LAYER metal1 ;
        RECT 2.6 6.3 3 6.7 ;
        RECT 0.6 3.4 6.4 3.7 ;
        RECT 6 3.3 6.4 3.7 ;
        RECT 2.6 3.4 3 3.8 ;
        RECT 2.1 2.3 2.5 2.7 ;
        RECT 2 2.7 2.4 3.7 ;
        RECT 0.6 3.3 1.4 3.7 ;
        RECT 2.7 6.7 3.1 7.1 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.4 4.2 1.8 4.6 ;
        RECT 3.4 4.3 3.8 4.7 ;
        RECT 1.4 4.3 3.8 4.6 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 2.6 ;
        RECT -0.2 -0.3 9.8 0.3 ;
        RECT 8.2 -0.3 8.6 2.5 ;
        RECT 5.4 -0.3 5.8 1.6 ;
        RECT 3.7 -0.3 4.2 1.6 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 5.5 1.4 10.3 ;
        RECT -0.2 9.7 9.8 10.3 ;
        RECT 8.2 5.4 8.6 10.3 ;
        RECT 5.4 7.4 5.8 10.3 ;
        RECT 3.8 7.4 4.2 10.3 ;
    END
  END vdd
  OBS
    LAYER metal2 ;
      RECT 0.2 2.6 0.6 5.4 ;
      RECT 1.8 1.6 2.2 5 ;
      RECT 1.8 1.6 2.1 7.4 ;
      RECT 1.8 5.4 2.2 7.4 ;
      RECT 6.6 1.6 7 5.7 ;
      RECT 6.6 1.6 6.9 7.4 ;
      RECT 6.6 6.1 7 7.4 ;
    LAYER metal1 ;
      RECT 0.2 0.6 0.6 3 ;
      RECT 1.8 7 2.2 7.7 ;
      RECT 1.8 7.4 2.8 7.7 ;
      RECT 2.4 7.4 2.8 9.4 ;
      RECT 2.4 0.6 2.8 1.6 ;
      RECT 1.8 1.3 2.8 1.6 ;
      RECT 1.8 1.3 2.2 2 ;
      RECT 1.8 5.7 4.5 6 ;
      RECT 1.8 5.7 2.2 6.1 ;
      RECT 4.1 5.7 4.5 6.1 ;
      RECT 4.6 0.6 5 1.6 ;
      RECT 4.6 0.6 4.9 2.2 ;
      RECT 3.5 1.9 4.9 2.2 ;
      RECT 3.5 1.9 3.9 2.3 ;
      RECT 3.5 6.7 3.9 7.1 ;
      RECT 4.9 6.7 5.3 7.1 ;
      RECT 3.5 6.8 5.3 7.1 ;
      RECT 4.6 6.8 4.9 9.4 ;
      RECT 4.6 7.4 5 9.4 ;
      RECT 6.6 7 7 7.4 ;
      RECT 6.7 7.4 7.3 9.4 ;
      RECT 0.2 4.9 2.5 5.2 ;
      RECT 2.1 5.1 5.7 5.4 ;
      RECT 5.4 5.1 5.7 6.1 ;
      RECT 5.4 5.7 7.3 6 ;
      RECT 5.4 5.7 5.9 6.1 ;
      RECT 6.9 5.7 7.3 6.1 ;
      RECT 0.2 4.9 0.6 9.4 ;
      RECT 6.7 0.6 7.3 1.6 ;
      RECT 6.6 1.3 7 2 ;
      RECT 6.6 4 7 4.4 ;
      RECT 6.6 4.1 8.5 4.4 ;
      RECT 8.1 4.1 8.5 4.5 ;
    LAYER via ;
      RECT 0.3 5.1 0.5 5.3 ;
      RECT 0.3 2.7 0.5 2.9 ;
      RECT 1.9 7.1 2.1 7.3 ;
      RECT 1.9 5.8 2.1 6 ;
      RECT 1.9 1.7 2.1 1.9 ;
      RECT 6.7 7.1 6.9 7.3 ;
      RECT 6.7 4.1 6.9 4.3 ;
      RECT 6.7 1.7 6.9 1.9 ;
  END
END DFFNEGX1

MACRO DFFPOSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFPOSX1 0 0 ;
  SIZE 9.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.3 4.7 7.7 5.1 ;
        RECT 9 0.6 9.4 9.4 ;
        RECT 7.3 4.8 9.4 5.1 ;
        RECT 7.5 2.8 9.4 3.1 ;
        RECT 7.5 2.7 7.9 3.1 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 0.6 3.3 1.4 3.7 ;
        RECT 6.7 6.1 7.4 6.5 ;
        RECT 6.7 5.3 7 6.5 ;
        RECT 5.8 5.3 7 5.6 ;
        RECT 5.8 3.4 6.1 5.6 ;
        RECT 5.5 3.3 5.9 3.7 ;
        RECT 0.6 3.4 6.1 3.7 ;
        RECT 2.7 1.9 3 3.7 ;
        RECT 2.6 1.9 3 2.3 ;
        RECT 2.1 3.4 2.5 3.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.3 4.2 1.7 4.6 ;
        RECT 3.4 4.3 3.8 4.7 ;
        RECT 1.3 4.3 3.8 4.6 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 2.6 ;
        RECT -0.2 -0.3 9.8 0.3 ;
        RECT 8.2 -0.3 8.6 2.5 ;
        RECT 5.4 -0.3 5.8 1.6 ;
        RECT 3.7 -0.3 4.2 1.6 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 5.5 1.4 10.3 ;
        RECT -0.2 9.7 9.8 10.3 ;
        RECT 8.2 5.4 8.6 10.3 ;
        RECT 5.4 7.4 5.8 10.3 ;
        RECT 3.8 7.4 4.2 10.3 ;
    END
  END vdd
  OBS
    LAYER metal2 ;
      RECT 0.2 2.6 0.6 5.4 ;
      RECT 1.8 1.6 2.2 7.4 ;
      RECT 6.6 1.6 7 7.4 ;
    LAYER metal1 ;
      RECT 0.2 0.6 0.6 3 ;
      RECT 1.8 7 2.2 7.7 ;
      RECT 1.8 7.4 2.8 7.7 ;
      RECT 2.4 7.4 2.8 9.4 ;
      RECT 2.4 0.6 2.8 1.6 ;
      RECT 1.8 1.3 2.8 1.6 ;
      RECT 1.8 1.3 2.2 2 ;
      RECT 1.8 5.7 4.5 6 ;
      RECT 1.8 5.7 2.2 6.1 ;
      RECT 4.1 5.7 4.5 6.1 ;
      RECT 4.6 0.6 5 1.6 ;
      RECT 4.6 0.6 4.9 2.2 ;
      RECT 3.5 1.9 4.9 2.2 ;
      RECT 3.5 1.9 3.9 2.3 ;
      RECT 3.5 6.7 3.9 7.1 ;
      RECT 4.9 6.7 5.3 7.1 ;
      RECT 3.5 6.8 5.3 7.1 ;
      RECT 4.6 6.8 4.9 9.4 ;
      RECT 4.6 7.4 5 9.4 ;
      RECT 0.2 5 3.1 5.2 ;
      RECT 0.2 4.9 3 5.2 ;
      RECT 2.7 5.1 5.1 5.4 ;
      RECT 4.8 5.1 5.1 6.3 ;
      RECT 5.5 5.9 5.9 6.3 ;
      RECT 4.8 6 5.9 6.3 ;
      RECT 0.2 4.9 0.6 9.4 ;
      RECT 6.6 7 7 7.4 ;
      RECT 6.7 7.4 7.3 9.4 ;
      RECT 6.7 0.6 7.3 1.6 ;
      RECT 6.6 1.3 7 2 ;
      RECT 6.6 4 7 4.4 ;
      RECT 6.6 4.1 8.5 4.4 ;
      RECT 8.1 4.1 8.5 4.5 ;
    LAYER via ;
      RECT 0.3 5.1 0.5 5.3 ;
      RECT 0.3 2.7 0.5 2.9 ;
      RECT 1.9 7.1 2.1 7.3 ;
      RECT 1.9 5.8 2.1 6 ;
      RECT 1.9 1.7 2.1 1.9 ;
      RECT 6.7 7.1 6.9 7.3 ;
      RECT 6.7 4.1 6.9 4.3 ;
      RECT 6.7 1.7 6.9 1.9 ;
  END
END DFFPOSX1

MACRO DFFSR
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSR 0 0 ;
  SIZE 17.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 16.2 0.6 16.6 2.9 ;
        RECT 16.3 2.5 16.7 5.5 ;
        RECT 16.2 5.1 16.6 9.4 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 8.2 2.3 9 2.7 ;
    END
  END CLK
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.9 4.4 1.3 4.8 ;
        RECT 0.9 4.5 12.6 4.8 ;
        RECT 12.2 4.2 12.6 4.8 ;
        RECT 3.4 4.3 3.8 4.8 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 5.1 2.2 5.7 ;
        RECT 1.8 5.1 15.3 5.4 ;
        RECT 14.9 5 15.3 5.4 ;
        RECT 3.5 5.1 3.9 5.5 ;
    END
  END S
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.6 2.9 7 3.7 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.8 -0.3 2.2 2.6 ;
        RECT -0.2 -0.3 17.8 0.3 ;
        RECT 17 -0.3 17.4 1.6 ;
        RECT 13.8 -0.3 14.2 2.6 ;
        RECT 8.2 -0.3 8.6 1.6 ;
        RECT 6.6 -0.3 7 1.6 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 7.4 0.6 10.3 ;
        RECT -0.2 9.7 17.8 10.3 ;
        RECT 17 7.4 17.4 10.3 ;
        RECT 15.4 7.4 15.8 10.3 ;
        RECT 13.8 7.4 14.2 10.3 ;
        RECT 12.2 7.4 12.6 10.3 ;
        RECT 8.2 7.4 8.6 10.3 ;
        RECT 6.6 7.4 7 10.3 ;
        RECT 3.4 7.4 3.8 10.3 ;
        RECT 1.8 7.4 2.2 10.3 ;
    END
  END vdd
  OBS
    LAYER metal2 ;
      RECT 4.2 1.6 4.6 8.4 ;
      RECT 5 1.6 5.4 8.4 ;
      RECT 5.8 1.6 6.2 7.4 ;
      RECT 7.4 1.6 7.8 7.4 ;
      RECT 9 1.6 9.4 7.4 ;
      RECT 9.8 1.6 10.2 8.4 ;
      RECT 10.6 1.6 11 8.4 ;
      RECT 11.4 1.6 11.8 8.4 ;
    LAYER metal1 ;
      RECT 3.4 0.6 3.8 2.6 ;
      RECT 2.5 2.2 3.8 2.6 ;
      RECT 2.5 2.2 2.9 3.3 ;
      RECT 1.4 2.9 2.9 3.3 ;
      RECT 4.2 8 4.6 9.4 ;
      RECT 0.2 3.6 4.6 4 ;
      RECT 0.2 0.6 0.6 7.1 ;
      RECT 0.2 6.8 1.2 7.1 ;
      RECT 0.9 6.8 1.2 7.7 ;
      RECT 1 7.4 1.4 9.4 ;
      RECT 4.2 0.6 4.6 2 ;
      RECT 5 8 5.4 9.4 ;
      RECT 2.7 5.8 5.4 6.1 ;
      RECT 5 5.7 5.4 6.1 ;
      RECT 2.3 6 3 6.4 ;
      RECT 5 0.6 5.4 2 ;
      RECT 5.8 7 6.2 9.4 ;
      RECT 5.8 0.6 6.2 2 ;
      RECT 7.4 7 7.8 9.4 ;
      RECT 6.5 6.3 7.8 6.7 ;
      RECT 5.5 2.3 7.8 2.6 ;
      RECT 7.4 2.3 7.8 2.7 ;
      RECT 5.5 2.3 5.9 4.2 ;
      RECT 4.9 3.8 5.9 4.2 ;
      RECT 7.4 0.6 7.8 2 ;
      RECT 9 6.3 9.4 9.4 ;
      RECT 7.8 3.8 9.4 4.2 ;
      RECT 9 0.6 9.4 2 ;
      RECT 7.4 3 7.8 3.4 ;
      RECT 7.4 3.1 9.6 3.4 ;
      RECT 9.2 3.1 9.6 3.5 ;
      RECT 9.8 8 10.2 9.4 ;
      RECT 5.9 5.7 10.2 6 ;
      RECT 9.8 5.7 10.2 6.1 ;
      RECT 1 6.1 1.8 6.5 ;
      RECT 1.5 6.1 1.8 7.1 ;
      RECT 3.3 6.4 6.2 6.7 ;
      RECT 5.9 5.7 6.2 6.7 ;
      RECT 1.5 6.7 3.6 7.1 ;
      RECT 2.6 6.7 3 9.4 ;
      RECT 9.8 0.6 10.2 2 ;
      RECT 10.6 8 11 9.4 ;
      RECT 10.5 2.3 11 2.7 ;
      RECT 10.6 2.3 11 4.1 ;
      RECT 10.6 0.6 11 2 ;
      RECT 11.4 8 11.8 9.4 ;
      RECT 11.4 0.6 11.8 2 ;
      RECT 10.6 6.7 12.7 7.1 ;
      RECT 13 6.3 14.3 6.7 ;
      RECT 13 6.3 13.4 9.4 ;
      RECT 12.2 0.6 12.6 2.6 ;
      RECT 12.2 2.2 13.4 2.6 ;
      RECT 13 2.2 13.4 3.2 ;
      RECT 13 2.9 13.9 3.2 ;
      RECT 13.5 2.9 13.9 4.2 ;
      RECT 13.5 3.8 15.4 4.2 ;
      RECT 15.4 0.6 15.8 3.5 ;
      RECT 15.7 3.2 16 4.8 ;
      RECT 11.4 5.7 15.9 6 ;
      RECT 11.4 5.7 11.8 6.1 ;
      RECT 15.6 4.5 15.9 7.1 ;
      RECT 14.6 6.8 15.9 7.1 ;
      RECT 14.6 6.8 15 9.4 ;
    LAYER via ;
      RECT 4.3 8.1 4.5 8.3 ;
      RECT 4.3 3.7 4.5 3.9 ;
      RECT 4.3 1.7 4.5 1.9 ;
      RECT 5.1 8.1 5.3 8.3 ;
      RECT 5.1 5.8 5.3 6 ;
      RECT 5.1 1.7 5.3 1.9 ;
      RECT 5.9 7.1 6.1 7.3 ;
      RECT 5.9 1.7 6.1 1.9 ;
      RECT 7.5 7.1 7.7 7.3 ;
      RECT 7.5 6.4 7.7 6.6 ;
      RECT 7.5 3.1 7.7 3.3 ;
      RECT 7.5 1.7 7.7 1.9 ;
      RECT 9.1 7.1 9.3 7.3 ;
      RECT 9.1 3.9 9.3 4.1 ;
      RECT 9.1 1.7 9.3 1.9 ;
      RECT 9.9 8.1 10.1 8.3 ;
      RECT 9.9 5.8 10.1 6 ;
      RECT 9.9 1.7 10.1 1.9 ;
      RECT 10.7 8.1 10.9 8.3 ;
      RECT 10.7 6.8 10.9 7 ;
      RECT 10.7 1.7 10.9 1.9 ;
      RECT 11.5 8.1 11.7 8.3 ;
      RECT 11.5 5.8 11.7 6 ;
      RECT 11.5 1.7 11.7 1.9 ;
  END
END DFFSR

MACRO FAX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FAX1 0 0 ;
  SIZE 12 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 11.4 0.6 11.8 1.6 ;
        RECT 11.4 7.4 11.8 9.4 ;
        RECT 11.5 0.6 11.8 9.4 ;
        RECT 11.4 3.3 11.8 3.7 ;
    END
  END YC
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.8 0.6 10.2 1.6 ;
        RECT 10.4 2.3 11 2.7 ;
        RECT 9.7 4.6 10.7 4.9 ;
        RECT 10.4 1.9 10.7 4.9 ;
        RECT 9.9 1.9 10.7 2.2 ;
        RECT 9.8 7.4 10.2 9.4 ;
        RECT 9.9 0.6 10.2 2.2 ;
        RECT 9.7 4.6 10 7.7 ;
    END
  END YS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3 3 1 3.3 ;
        RECT 8.9 3.4 9.3 3.8 ;
        RECT 8.9 2.8 9.2 3.8 ;
        RECT 3.7 2.8 9.2 3.1 ;
        RECT 0.3 3 4.1 3.2 ;
        RECT 0.6 2.9 9.2 3.1 ;
        RECT 0.2 3.3 0.6 3.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.1 3.6 1.4 4.7 ;
        RECT 8 3.4 8.4 3.8 ;
        RECT 4.7 3.4 8.4 3.7 ;
        RECT 1.1 3.6 5.1 3.8 ;
        RECT 1.4 3.5 8.4 3.7 ;
        RECT 2.9 3.5 3.3 3.9 ;
        RECT 1.1 3.6 1.8 3.9 ;
        RECT 1 4.3 1.4 4.7 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 4.3 2.6 4.7 ;
        RECT 7.2 4 7.6 4.4 ;
        RECT 5.2 4.1 7.6 4.4 ;
        RECT 1.8 4.3 5.9 4.5 ;
        RECT 1.8 4.3 5.5 4.6 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 2 ;
        RECT -0.2 -0.3 12.2 0.3 ;
        RECT 10.6 -0.3 11 1.6 ;
        RECT 9 -0.3 9.4 2.5 ;
        RECT 5.5 -0.3 5.9 1.9 ;
        RECT 3.9 -0.3 4.3 2.4 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 6 1.4 10.3 ;
        RECT -0.2 9.7 12.2 10.3 ;
        RECT 10.6 7.4 11 10.3 ;
        RECT 9 4.6 9.4 10.3 ;
        RECT 5.5 6.4 5.9 10.3 ;
        RECT 3.9 5.4 4.3 10.3 ;
    END
  END vdd
  OBS
    LAYER metal2 ;
      RECT 7.2 2.1 7.6 2.5 ;
      RECT 7.3 3.9 10.1 4.2 ;
      RECT 9.7 3.9 10.1 4.3 ;
      RECT 7.3 2.1 7.6 5.1 ;
      RECT 7.2 4.7 7.6 5.1 ;
      RECT 2.6 2.2 3 2.6 ;
      RECT 6 4.8 6.4 5.7 ;
      RECT 10.4 5.3 10.8 5.7 ;
      RECT 2.6 5.4 10.8 5.7 ;
      RECT 2.7 2.2 3 5.8 ;
      RECT 2.6 5.4 3 5.8 ;
    LAYER metal1 ;
      RECT 0.2 5.4 2.2 5.7 ;
      RECT 0.2 5.4 0.6 9.4 ;
      RECT 1.8 5.4 2.2 9.4 ;
      RECT 0.2 0.6 0.6 2.6 ;
      RECT 1.8 0.6 2.2 2.6 ;
      RECT 0.2 2.3 2.2 2.6 ;
      RECT 2.6 5.4 3 9.4 ;
      RECT 2.6 0.6 3 2.6 ;
      RECT 4.7 5.8 6.7 6.1 ;
      RECT 4.7 5.4 5.1 9.4 ;
      RECT 6.3 5.8 6.7 9.4 ;
      RECT 4.7 0.6 5.1 2.5 ;
      RECT 6.3 0.6 6.7 2.5 ;
      RECT 4.7 2.2 6.7 2.5 ;
      RECT 6.4 4.7 6.8 5.1 ;
      RECT 6 4.8 6.4 5.2 ;
      RECT 7.2 4.7 7.6 9.4 ;
      RECT 7.1 5.1 7.6 9.4 ;
      RECT 7.1 0.6 7.6 2.1 ;
      RECT 7.2 0.6 7.6 2.5 ;
      RECT 9.7 3.5 10.1 4.3 ;
      RECT 10.4 5.3 11.2 5.7 ;
    LAYER via ;
      RECT 2.7 5.5 2.9 5.7 ;
      RECT 2.7 2.3 2.9 2.5 ;
      RECT 6.1 4.9 6.3 5.1 ;
      RECT 7.3 4.8 7.5 5 ;
      RECT 7.3 2.2 7.5 2.4 ;
      RECT 9.8 4 10 4.2 ;
      RECT 10.5 5.4 10.7 5.6 ;
  END
END FAX1

MACRO FILL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL 0 0 ;
  SIZE 0.8 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.2 -0.3 1 0.3 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.2 9.7 1 10.3 ;
    END
  END vdd
END FILL

MACRO HAX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HAX1 0 0 ;
  SIZE 8 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 2.3 1.6 3 2 ;
        RECT 2.6 4.2 3 4.6 ;
        RECT 2.7 1.6 3 4.6 ;
      LAYER via ;
        RECT 2.4 1.7 2.6 1.9 ;
        RECT 2.7 4.3 2.9 4.5 ;
      LAYER metal1 ;
        RECT 2.3 0.6 2.7 2 ;
        RECT 2.6 4.2 3 9.4 ;
    END
  END YC
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.6 5.3 7 5.7 ;
        RECT 7.1 7.4 7.5 9.4 ;
        RECT 7.2 6.8 7.5 9.4 ;
        RECT 6.7 2 7.5 2.3 ;
        RECT 7.2 0.6 7.5 2.3 ;
        RECT 6.7 6.8 7.5 7.1 ;
        RECT 7.1 0.6 7.5 1.6 ;
        RECT 6.7 2 7 7.1 ;
    END
  END YS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3 0.6 3.7 ;
        RECT 5 3.3 5.4 3.7 ;
        RECT 4.2 3.3 5.4 3.6 ;
        RECT 0.2 3 4.5 3.3 ;
        RECT 0.4 2.9 0.8 3.3 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.1 4 1.5 4.3 ;
        RECT 4.2 3.9 4.6 4.3 ;
        RECT 3.6 3.9 4.6 4.2 ;
        RECT 1.2 3.6 3.9 3.9 ;
        RECT 1.2 3.6 1.6 4 ;
        RECT 1 4.3 1.4 4.7 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 2.6 ;
        RECT -0.2 -0.3 8.2 0.3 ;
        RECT 6.3 -0.3 6.7 1.6 ;
        RECT 3.1 -0.3 3.5 2.5 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 7.6 1.4 10.3 ;
        RECT -0.2 9.7 8.2 10.3 ;
        RECT 6.3 7.4 6.7 10.3 ;
        RECT 5.5 5.4 5.9 10.3 ;
        RECT 3.4 7.4 3.8 10.3 ;
    END
  END vdd
  OBS
    LAYER metal2 ;
      RECT 1.9 2.3 2.3 2.7 ;
      RECT 1.9 2.3 2.2 4.6 ;
      RECT 1.9 4.2 2.3 4.6 ;
    LAYER metal1 ;
      RECT 1.9 4.2 2.3 4.6 ;
      RECT 0.3 7 2.2 7.3 ;
      RECT 0.3 7 0.6 9.4 ;
      RECT 0.2 7.4 0.6 9.4 ;
      RECT 1.9 4.2 2.2 9.4 ;
      RECT 1.8 7 2.2 9.4 ;
      RECT 1.5 0.6 1.9 2.6 ;
      RECT 1.9 2.3 2.8 2.7 ;
      RECT 3.9 0.6 5.9 0.9 ;
      RECT 5.5 0.6 5.9 2.4 ;
      RECT 3.9 0.6 4.3 2.6 ;
      RECT 4.7 1.2 5.1 2.6 ;
      RECT 4.8 1.2 5.1 3 ;
      RECT 4.8 2.7 6.3 3 ;
      RECT 5.7 2.7 6.3 3.1 ;
      RECT 5.7 2.7 6 5.1 ;
      RECT 4.3 4.8 6 5.1 ;
      RECT 4.3 4.8 4.6 9.4 ;
      RECT 4.2 5.4 4.6 9.4 ;
    LAYER via ;
      RECT 2 4.3 2.2 4.5 ;
      RECT 2 2.4 2.2 2.6 ;
  END
END HAX1

MACRO INVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1 0 0 ;
  SIZE 1.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 1.9 0.6 2.7 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 1.6 ;
        RECT -0.2 -0.3 1.8 0.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 0.6 1.4 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 7.4 0.6 10.3 ;
        RECT -0.2 9.7 1.8 10.3 ;
    END
  END vdd
END INVX1

MACRO INVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2 0 0 ;
  SIZE 1.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 2.9 0.6 3.7 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 2.6 ;
        RECT -0.2 -0.3 1.8 0.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 0.6 1.4 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 1.8 10.3 ;
    END
  END vdd
END INVX2

MACRO INVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX4 0 0 ;
  SIZE 2.4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 2.9 0.6 3.7 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 2.6 ;
        RECT -0.2 -0.3 2.6 0.3 ;
        RECT 1.8 -0.3 2.2 2.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 0.6 1.4 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 2.6 10.3 ;
        RECT 1.8 5.4 2.2 10.3 ;
    END
  END vdd
END INVX4

MACRO INVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX8 0 0 ;
  SIZE 4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 2.9 0.6 3.7 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 2.6 ;
        RECT -0.2 -0.3 4.2 0.3 ;
        RECT 3.4 -0.3 3.8 2.6 ;
        RECT 1.8 -0.3 2.2 2.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 0.6 1.4 3.3 ;
        RECT 2.6 0.6 3 9.4 ;
        RECT 1 4.7 3 5.1 ;
        RECT 1 2.9 3 3.3 ;
        RECT 1 4.7 1.4 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 4.2 10.3 ;
        RECT 3.4 5.4 3.8 10.3 ;
        RECT 1.8 5.4 2.2 10.3 ;
    END
  END vdd
END INVX8

MACRO LATCH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATCH 0 0 ;
  SIZE 5.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.7 3.8 5.4 4.2 ;
        RECT 5 0.6 5.4 9.4 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 0.6 3.3 1.4 3.7 ;
        RECT 2.9 3.3 3.3 4.1 ;
        RECT 0.6 3.3 3.3 3.6 ;
        RECT 2.2 2.3 2.6 3.6 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.3 4.7 2.2 5.1 ;
        RECT 1.8 4.7 2.2 5.7 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 2.6 ;
        RECT -0.2 -0.3 5.8 0.3 ;
        RECT 4.2 -0.3 4.6 2.6 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 5.4 1.4 10.3 ;
        RECT -0.2 9.7 5.8 10.3 ;
        RECT 4.2 5.4 4.6 10.3 ;
    END
  END vdd
  OBS
    LAYER metal2 ;
      RECT 0.2 2.6 0.6 5.4 ;
      RECT 2.6 1.6 3 7.4 ;
    LAYER metal1 ;
      RECT 0.2 4.9 0.6 9.4 ;
      RECT 0.2 0.6 0.6 3 ;
      RECT 0.2 4 2.5 4.3 ;
      RECT 0.2 4 0.6 4.4 ;
      RECT 2.1 4 2.5 4.4 ;
      RECT 2.6 7 3 9.4 ;
      RECT 2.5 7.4 3.1 9.4 ;
      RECT 2.5 0.6 3.1 1.6 ;
      RECT 2.6 0.6 3 2 ;
      RECT 2.6 4.7 4.7 5.1 ;
    LAYER via ;
      RECT 0.3 5.1 0.5 5.3 ;
      RECT 0.3 4.1 0.5 4.3 ;
      RECT 0.3 2.7 0.5 2.9 ;
      RECT 2.7 7.1 2.9 7.3 ;
      RECT 2.7 4.8 2.9 5 ;
      RECT 2.7 1.7 2.9 1.9 ;
  END
END LATCH

MACRO MUX2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X1 0 0 ;
  SIZE 4.8 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.4 4.3 3.8 5.1 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 3.9 1.4 4.7 ;
    END
  END B
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.9 0.6 4.7 ;
    END
  END S
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 2.8 ;
        RECT -0.2 -0.3 5 0.3 ;
        RECT 3.6 -0.3 4 3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.3 1 2.7 2.8 ;
        RECT 2.8 3.3 3.8 3.7 ;
        RECT 2.3 5.6 3.1 5.9 ;
        RECT 2.8 2.5 3.1 5.9 ;
        RECT 2.7 2.5 3.1 3 ;
        RECT 2.3 5.6 2.7 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 5.6 1.4 10.3 ;
        RECT -0.2 9.7 5 10.3 ;
        RECT 3.6 5.4 4 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.2 1 0.6 2 ;
      RECT 0.2 1 0.5 3.4 ;
      RECT 0.2 3.1 2.3 3.4 ;
      RECT 1.8 3.1 2.3 4 ;
      RECT 1.8 3.6 2.5 4 ;
      RECT 1.8 3.1 2.1 5.3 ;
      RECT 0.2 5 2.1 5.3 ;
      RECT 0.2 5 0.5 9 ;
      RECT 0.2 7 0.6 9 ;
  END
END MUX2X1

MACRO NAND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1 0 0 ;
  SIZE 2.4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 2.9 0.6 3.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 5.3 2.2 6.1 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 2.6 ;
        RECT -0.2 -0.3 2.6 0.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 2.3 1.4 9.4 ;
        RECT 1 2.3 1.9 2.6 ;
        RECT 1.5 0.6 1.9 2.6 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 7.4 0.6 10.3 ;
        RECT -0.2 9.7 2.6 10.3 ;
        RECT 1.8 7.4 2.2 10.3 ;
    END
  END vdd
END NAND2X1

MACRO NAND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X1 0 0 ;
  SIZE 3.2 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 4.9 0.6 5.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 4.3 1.8 4.7 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 5.9 2.2 6.7 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 3.6 ;
        RECT -0.2 -0.3 3.4 0.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.1 7 1.4 9.4 ;
        RECT 2.6 7.4 3 9.4 ;
        RECT 2.6 5.3 3 5.7 ;
        RECT 2.6 3.4 2.9 9.4 ;
        RECT 1.1 7 2.9 7.3 ;
        RECT 2.1 3.4 2.9 3.7 ;
        RECT 2 0.6 2.4 3.6 ;
        RECT 1 7.4 1.4 9.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 7.4 0.6 10.3 ;
        RECT -0.2 9.7 3.4 10.3 ;
        RECT 1.8 7.6 2.2 10.3 ;
    END
  END vdd
END NAND3X1

MACRO NOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X1 0 0 ;
  SIZE 2.4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 1.9 0.6 2.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 4.3 2.2 5.1 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 1.6 ;
        RECT -0.2 -0.3 2.6 0.3 ;
        RECT 1.8 -0.3 2.2 1.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 0.6 1.4 1.6 ;
        RECT 1.5 5.4 1.9 9.4 ;
        RECT 1 5.4 1.9 5.8 ;
        RECT 1.1 0.6 1.4 5.8 ;
        RECT 1 3.3 1.4 3.7 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 2.6 10.3 ;
    END
  END vdd
END NOR2X1

MACRO NOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X1 0 0 ;
  SIZE 6.4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 2.3 1.9 2.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 3.3 2.6 3.7 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6 4.3 3.4 4.7 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 1.6 ;
        RECT -0.2 -0.3 6.6 0.3 ;
        RECT 2.6 -0.3 3 1.4 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 0.6 2.2 1.6 ;
        RECT 5 6 5.4 8.8 ;
        RECT 5 5.3 5.4 5.7 ;
        RECT 5 5.3 5.3 8.8 ;
        RECT 3.7 5.3 5.4 5.6 ;
        RECT 3.7 1.6 4 5.6 ;
        RECT 3.4 0.6 3.8 2 ;
        RECT 2 1.7 4 2 ;
        RECT 2 1.3 2.3 2 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 6.4 1.4 10.3 ;
        RECT -0.2 9.7 6.6 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.3 5.8 2.1 6.1 ;
      RECT 1.8 5.8 2.1 9.4 ;
      RECT 1.8 6.4 2.2 9.4 ;
      RECT 0.3 5.8 0.6 9.4 ;
      RECT 0.2 6.4 0.6 9.4 ;
      RECT 3.4 6.5 3.8 9.4 ;
      RECT 1.8 9.1 3.8 9.4 ;
      RECT 2.7 5.9 4.5 6.2 ;
      RECT 2.7 5.9 3 8.8 ;
      RECT 2.6 6.4 3 8.8 ;
      RECT 4.2 6 4.6 9 ;
      RECT 5.8 6 6.2 9 ;
      RECT 4.3 6 4.6 9.4 ;
      RECT 5.8 6 6.1 9.4 ;
      RECT 4.3 9.1 6.1 9.4 ;
  END
END NOR3X1

MACRO OAI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X1 0 0 ;
  SIZE 3.2 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.3 0.6 3.7 ;
        RECT 0.6 3.1 1 3.6 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 3.9 1.4 4.7 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.3 5.4 2.6 6.7 ;
        RECT 2.6 5.3 3 5.7 ;
        RECT 2.2 6.3 2.6 6.7 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 2.2 ;
        RECT -0.2 -0.3 3.4 0.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.5 5.4 1.9 9.4 ;
        RECT 1.7 3.3 3 3.7 ;
        RECT 2.6 0.6 3 2.6 ;
        RECT 2.6 0.6 2.9 3.7 ;
        RECT 1.7 3.3 2 5.7 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 3.4 10.3 ;
        RECT 2.3 7.4 2.7 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.2 0.6 0.6 2.6 ;
      RECT 1.8 0.6 2.2 2.6 ;
      RECT 0.3 2.5 2.1 2.8 ;
  END
END OAI21X1

MACRO OAI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X1 0 0 ;
  SIZE 4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.3 0.6 3.7 ;
        RECT 0.6 3.1 1 3.6 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 3.9 1.4 4.7 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.4 3.3 3.8 4.1 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6 3.9 3 4.7 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 -0.3 1.4 2.2 ;
        RECT -0.2 -0.3 4.2 0.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 3.3 2.1 9.4 ;
        RECT 1.8 3.3 3 3.6 ;
        RECT 2.7 1.2 3 3.6 ;
        RECT 2.6 1.2 3 2.6 ;
        RECT 1.5 5.4 2.5 9.4 ;
        RECT 1.8 3.3 2.2 3.7 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 4.2 10.3 ;
        RECT 3.4 5.4 3.8 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 1.8 0.6 3.8 0.9 ;
      RECT 0.2 0.6 0.6 2.6 ;
      RECT 1.8 0.6 2.2 2.6 ;
      RECT 3.4 0.6 3.8 2.6 ;
      RECT 0.3 2.5 2.1 2.8 ;
  END
END OAI22X1

MACRO OR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X1 0 0 ;
  SIZE 3.2 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 1.9 0.6 2.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 3.3 1.4 3.7 ;
        RECT 1.1 2.9 1.8 3.3 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 1.6 ;
        RECT -0.2 -0.3 3.4 0.3 ;
        RECT 1.8 -0.3 2.2 1.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6 0.6 3 1.6 ;
        RECT 2.7 0.6 3 7.4 ;
        RECT 2.3 7.4 2.7 9.4 ;
        RECT 2.4 7.1 3 7.4 ;
        RECT 2.6 4.3 3 4.7 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.5 5.4 1.9 10.3 ;
        RECT -0.2 9.7 3.4 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 1 0.6 1.4 1.6 ;
      RECT 1.1 0.6 1.4 2.4 ;
      RECT 1.1 2.1 2.4 2.4 ;
      RECT 2.1 2.1 2.4 3.9 ;
      RECT 1.9 3.6 2.2 5.1 ;
      RECT 1.9 4.7 2.3 5.1 ;
      RECT 0.2 4.8 2.3 5.1 ;
      RECT 0.2 4.8 0.6 9.4 ;
  END
END OR2X1

MACRO OR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X2 0 0 ;
  SIZE 3.2 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 1.9 0.6 2.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1 3.3 1.5 3.7 ;
        RECT 1.2 3.7 1.6 4.1 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 1.6 ;
        RECT -0.2 -0.3 3.4 0.3 ;
        RECT 1.8 -0.3 2.2 2.4 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6 0.6 3 2.6 ;
        RECT 2.7 0.6 3 5.7 ;
        RECT 2.3 5.4 2.7 9.4 ;
        RECT 2.6 4.3 3 4.7 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.5 5.4 1.9 10.3 ;
        RECT -0.2 9.7 3.4 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 1 0.6 1.4 1.6 ;
      RECT 1.1 0.6 1.4 3 ;
      RECT 1.1 2.7 2.3 3 ;
      RECT 1.9 4.5 2.3 4.9 ;
      RECT 2 2.7 2.3 4.9 ;
      RECT 0.2 4.8 2.2 5.1 ;
      RECT 0.2 4.8 0.6 9.4 ;
  END
END OR2X2

MACRO TBUFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX1 0 0 ;
  SIZE 4 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 3.3 3.8 3.7 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 6.3 1 6.7 ;
    END
  END EN
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 1.6 ;
        RECT -0.2 -0.3 4.2 0.3 ;
        RECT 3.2 -0.3 3.6 2.6 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.9 0.6 2.3 2.6 ;
        RECT 1.9 5.4 2.3 9.4 ;
        RECT 2 0.6 2.3 9.4 ;
        RECT 1.8 4.3 2.3 4.7 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 7.4 0.6 10.3 ;
        RECT -0.2 9.7 4.2 10.3 ;
        RECT 3.2 5.4 3.6 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 1 0.6 1.4 1.6 ;
      RECT 1.3 3.3 1.7 3.7 ;
      RECT 1.3 1.2 1.6 4 ;
      RECT 1.2 3.7 1.5 5.3 ;
      RECT 1.3 5 1.6 7.7 ;
      RECT 1 7.4 1.4 9.4 ;
  END
END TBUFX1

MACRO TBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX2 0 0 ;
  SIZE 5.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.5 3.3 5.4 3.7 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 2.9 0.5 5.1 ;
        RECT 0.2 2.9 0.7 3.3 ;
        RECT 0.2 4.3 0.6 5.1 ;
    END
  END EN
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 -0.3 0.6 2.6 ;
        RECT -0.2 -0.3 5.8 0.3 ;
        RECT 4.2 -0.3 4.6 2.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6 1.2 2.9 8.8 ;
        RECT 2.6 5.4 3 8.8 ;
        RECT 2.6 4.3 3 4.7 ;
        RECT 2.6 1.2 3 2.6 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2 5.4 0.6 10.3 ;
        RECT -0.2 9.7 5.8 10.3 ;
        RECT 4.2 6.1 4.6 10.3 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 1 0.6 1.4 2.6 ;
      RECT 1 4.1 1.4 4.5 ;
      RECT 1 0.6 1.3 9.4 ;
      RECT 1 5.4 1.4 9.4 ;
      RECT 3.4 5.4 5.4 5.8 ;
      RECT 1.8 5.4 2.2 9.4 ;
      RECT 3.4 5.4 3.8 9.4 ;
      RECT 1.8 9.1 3.8 9.4 ;
      RECT 5 5.4 5.4 9.4 ;
      RECT 1.8 0.6 3.8 0.9 ;
      RECT 5 0.6 5.4 2.3 ;
      RECT 3.4 0.6 3.8 2.9 ;
      RECT 1.8 0.6 2.2 2.6 ;
      RECT 5.1 0.6 5.4 2.9 ;
      RECT 3.4 2.6 5.4 2.9 ;
  END
END TBUFX2

MACRO XNOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X1 0 0 ;
  SIZE 5.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 1.8 2.7 2.2 3.1 ;
        RECT 3.5 2.7 3.9 3.1 ;
        RECT 1.8 2.7 3.9 3 ;
      LAYER via ;
        RECT 1.9 2.8 2.1 3 ;
        RECT 3.6 2.8 3.8 3 ;
      LAYER metal1 ;
        RECT 0.2 3.3 1 3.7 ;
        RECT 3.6 3.3 4 3.7 ;
        RECT 3.6 2.7 3.9 3.7 ;
        RECT 3.5 2.7 3.9 3.1 ;
        RECT 1.8 2.7 2.6 3.1 ;
        RECT 0.2 3.3 1.9 3.6 ;
        RECT 1.6 2.8 1.9 3.6 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.6 3.3 5.4 3.7 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.1 -0.3 1.5 2.3 ;
        RECT -0.2 -0.3 5.8 0.3 ;
        RECT 4.1 -0.3 4.6 2.3 ;
        RECT 1 0.6 1.5 2.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.4 0.6 3.2 2.4 ;
        RECT 3.1 4.3 3.8 4.7 ;
        RECT 3.1 4.1 3.4 5.7 ;
        RECT 2.4 5.4 3.2 9.4 ;
        RECT 2.9 0.6 3.2 4.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 6.1 1.5 9.4 ;
        RECT -0.2 9.7 5.8 10.3 ;
        RECT 4.1 6.1 4.6 10.3 ;
        RECT 1.1 6.1 1.5 10.3 ;
    END
  END vdd
  OBS
    LAYER metal2 ;
      RECT 0.9 2.6 1.3 3 ;
      RECT 0.9 2.6 1.2 5.8 ;
      RECT 0.9 5.4 1.3 5.8 ;
      RECT 4.2 2.6 4.6 3 ;
      RECT 2.2 3.4 4.6 3.7 ;
      RECT 2.2 3.4 2.6 3.8 ;
      RECT 4.3 2.6 4.6 5.8 ;
      RECT 4.2 5.4 4.6 5.8 ;
    LAYER metal1 ;
      RECT 0.2 0.6 0.6 2.9 ;
      RECT 0.2 2.6 1.3 2.9 ;
      RECT 0.9 2.6 1.3 3 ;
      RECT 2.2 3.4 2.6 3.8 ;
      RECT 2.2 3.4 2.5 4.4 ;
      RECT 1.2 4.1 2.5 4.4 ;
      RECT 1.2 4.1 1.6 4.5 ;
      RECT 2.3 4.7 2.7 5.1 ;
      RECT 1 4.8 2.7 5.1 ;
      RECT 0.2 5.4 1.3 5.7 ;
      RECT 1 4.8 1.3 5.8 ;
      RECT 0.9 5.4 1.3 5.8 ;
      RECT 0.2 5.4 0.6 9.4 ;
      RECT 4.2 5.4 5.4 5.7 ;
      RECT 4.2 5.4 4.6 5.8 ;
      RECT 5 5.4 5.4 9.4 ;
      RECT 5 0.6 5.4 2.9 ;
      RECT 4.2 2.6 5.4 2.9 ;
      RECT 4.2 2.6 4.6 3 ;
    LAYER via ;
      RECT 1 5.5 1.2 5.7 ;
      RECT 1 2.7 1.2 2.9 ;
      RECT 2.3 3.5 2.5 3.7 ;
      RECT 4.3 5.5 4.5 5.7 ;
      RECT 4.3 2.7 4.5 2.9 ;
  END
END XNOR2X1

MACRO XOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X1 0 0 ;
  SIZE 5.6 BY 10 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 3.3 1 3.7 ;
        RECT 2 3.5 2.4 3.9 ;
        RECT 1 3.5 2.4 3.8 ;
        RECT 0.2 3.4 1.3 3.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.6 3.3 5.4 3.7 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.1 -0.3 1.5 2.3 ;
        RECT -0.2 -0.3 5.8 0.3 ;
        RECT 4.1 -0.3 4.6 2.3 ;
        RECT 1 0.6 1.5 2.3 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6 4.3 3 4.7 ;
        RECT 2.4 5.4 3.2 9.4 ;
        RECT 2.9 0.6 3.2 3.7 ;
        RECT 2.7 3.4 3 9.4 ;
        RECT 2.4 0.6 3.2 2.4 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1 6.1 1.5 9.4 ;
        RECT -0.2 9.7 5.8 10.3 ;
        RECT 4.1 6.1 4.6 10.3 ;
        RECT 1.1 6.1 1.5 10.3 ;
    END
  END vdd
  OBS
    LAYER metal2 ;
      RECT 1.1 2.6 1.5 3 ;
      RECT 1.1 2.7 3.9 3 ;
      RECT 1.8 2.7 2.2 3.1 ;
      RECT 3.5 2.7 3.9 3.1 ;
      RECT 1.1 2.6 1.4 5.8 ;
      RECT 1.1 5.4 1.5 5.8 ;
      RECT 4.2 2.6 4.6 3 ;
      RECT 1.8 3.4 4.6 3.7 ;
      RECT 1.8 3.4 2.1 4.8 ;
      RECT 1.7 4.4 2.1 4.8 ;
      RECT 4.3 2.6 4.6 5.8 ;
      RECT 4.2 5.4 4.6 5.8 ;
    LAYER metal1 ;
      RECT 0.2 5.4 1.5 5.7 ;
      RECT 1.1 5.4 1.5 5.8 ;
      RECT 0.2 5.4 0.6 9.4 ;
      RECT 0.2 0.6 0.6 2.9 ;
      RECT 0.2 2.6 1.5 2.9 ;
      RECT 1.1 2.6 1.5 3 ;
      RECT 1.3 4.3 1.7 4.7 ;
      RECT 1.7 4.4 2.1 4.8 ;
      RECT 1.8 2.7 2.6 3.1 ;
      RECT 3.5 2.7 3.9 3.1 ;
      RECT 3.6 2.7 3.9 3.7 ;
      RECT 3.6 3.3 4 3.7 ;
      RECT 4.2 5.4 5.4 5.7 ;
      RECT 4.2 5.4 4.6 5.8 ;
      RECT 5 5.4 5.4 9.4 ;
      RECT 5 0.6 5.4 2.9 ;
      RECT 4.2 2.6 5.4 2.9 ;
      RECT 4.2 2.6 4.6 3 ;
    LAYER via ;
      RECT 1.2 5.5 1.4 5.7 ;
      RECT 1.2 2.7 1.4 2.9 ;
      RECT 1.8 4.5 2 4.7 ;
      RECT 1.9 2.8 2.1 3 ;
      RECT 3.6 2.8 3.8 3 ;
      RECT 4.3 5.5 4.5 5.7 ;
      RECT 4.3 2.7 4.5 2.9 ;
  END
END XOR2X1

END LIBRARY
