VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.05 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER nactive
  TYPE MASTERSLICE ;
END nactive

LAYER pactive
  TYPE MASTERSLICE ;
END pactive

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER cc
  TYPE CUT ;
  SPACING 0.45 ;
END cc

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1 ;
  WIDTH 0.3 ;
  SPACING 0.3 ;
  RESISTANCE RPERSQ 0.08 ;
  CAPACITANCE CPERSQDIST 3.8e-05 ;
  EDGECAPACITANCE 8e-05 ;
END metal1

LAYER via
  TYPE CUT ;
  SPACING 0.3 ;
END via

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.8 ;
  WIDTH 0.3 ;
  SPACING 0.3 ;
  RESISTANCE RPERSQ 0.08 ;
  CAPACITANCE CPERSQDIST 1.9e-05 ;
  EDGECAPACITANCE 6e-05 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.3 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1 ;
  WIDTH 0.3 ;
  SPACING 0.3 ;
  RESISTANCE RPERSQ 0.08 ;
  CAPACITANCE CPERSQDIST 1.3e-05 ;
  EDGECAPACITANCE 5.4e-05 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.4 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.8 ;
  WIDTH 0.3 ;
  SPACING 0.3 ;
  RESISTANCE RPERSQ 0.07 ;
  CAPACITANCE CPERSQDIST 8e-06 ;
  EDGECAPACITANCE 4.1e-05 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.3 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1 ;
  WIDTH 0.3 ;
  SPACING 0.3 ;
  RESISTANCE RPERSQ 0.07 ;
  CAPACITANCE CPERSQDIST 8e-06 ;
  EDGECAPACITANCE 2.4e-05 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.4 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.6 ;
  WIDTH 0.5 ;
  SPACING 0.5 ;
  RESISTANCE RPERSQ 0.03 ;
  CAPACITANCE CPERSQDIST 3e-06 ;
  EDGECAPACITANCE 2e-05 ;
END metal6

VIARULE viagen21 GENERATE
  LAYER metal1 ;
    WIDTH 0.3 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER metal2 ;
    WIDTH 0.3 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER via ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.5 BY 0.5 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal2 ;
    WIDTH 0.3 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER metal3 ;
    WIDTH 0.3 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.5 BY 0.5 ;
END viagen32

VIARULE viagen43 GENERATE
  LAYER metal3 ;
    WIDTH 0.3 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER metal4 ;
    WIDTH 0.3 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.6 BY 0.6 ;
END viagen43

VIARULE viagen54 GENERATE
  LAYER metal4 ;
    WIDTH 0.3 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER metal5 ;
    WIDTH 0.3 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER via4 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.5 BY 0.5 ;
END viagen54

VIARULE viagen65 GENERATE
  LAYER metal5 ;
    WIDTH 0.5 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER metal6 ;
    WIDTH 0.5 TO 60 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER via5 ;
    RECT -0.15 -0.15 0.15 0.15 ;
    SPACING 0.7 BY 0.7 ;
END viagen65

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal2 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M3_M2

VIA M4_M3 DEFAULT
  LAYER metal3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal4 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M4_M3

VIA M5_M4 DEFAULT
  LAYER metal4 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via4 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal5 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M5_M4

VIA M6_M5 DEFAULT
  LAYER metal5 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER via5 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER metal6 ;
    RECT -0.25 -0.25 0.25 0.25 ;
END M6_M5

SITE core
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.8 BY 10 ;
END core

END LIBRARY
